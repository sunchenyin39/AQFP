*AQFP_RAM_CELL

Iwb     0       wb          pwl(0 0 5p 1410u)
Iy      0       y           pwl(0 0 310p 0 320p 40u 380p 40u 390p 0 1110p 0 1120p -40u 1180p -40u 1190p 0)
Ix      0       x           pwl(0 0 310p 0 320p 40u 380p 40u 390p 0 660p 0 670p -40u 730p -40u 740p 0 1110p 0 1120p -40u 1180p -40u 1190p 0 1460p 0 1470p -40u 1530p -40u 1540p 0)
Id      0       d           pwl(0 0 10p 50u 320p 50u 330p 140u 390p 140u 400p 50u 1120p 50u 1130p -40u 1190p -40u 1200p 50u)
Iclk    0       clk         pwl(0 0 100p 0 110p 1.2m 190p 1.2m 200p 0 300p 0 310p 1.2m 390p 1.2m 400p 0 500p 0 510p 1.2m 590p 1.2m 600p 0 700p 0 710p 1.2m 790p 1.2m 800p 0 900p 0 910p 1.2m 990p 1.2m 1000p 0 1100p 0 1110p 1.2m 1190p 1.2m 1200p 0 1300p 0 1310p 1.2m 1390p 1.2m 1400p 0 1500p 0 1510p 1.2m 1590p 1.2m 1600p 0)
Irb     0       rb          pwl(0 0 5p 50u)
X1      x y d clk q wb rb   AQFP_RAM_CELL
Lout    q       0           6.8p

.subckt AQFP_RAM_CELL x y d clk q wb rb
.model jjmod jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
B1      1       0       jjmod       area=0.5
B2      2       0       jjmod       area=0.5
Lw1     1       3       1.39p
Lw2     3       2       1.42p
Lp1     3       4       0.256p
Lin1    4       0       9.04p
Lin2    4       0       8.41p

Lwb     wb      0       12.6p
Kw1     Lwb     Lw1     -0.168
Kw2     Lwb     Lw2     -0.18

Ly      y       0       16.8p
Ky      Ly      Lin1    -0.301

Lx      x       0       16.1p
Kxw     Lx      Lin1    -0.157

Ld      d       0       13.1p
Kd      Ld      Lin2    -0.182

B3      9       0       jjmod       area=0.5
B4      10      0       jjmod       area=0.5
Lr1     9       11      1.36p   
Lr2     11      10      1.38p
Lqr     11      q       8.28p
Lp2     11      12      1.19p
Lin3    12      0       30.8p
Lin4    12      0       22.2p
Lclk    clk      0      14.2p
Kr1     Lclk    Lr1     -0.166
Kr2     Lclk    Lr2     -0.168

Lrb     rb      0       19.9p
Krb     Lrb     Lin4    -0.179
Kwr     Lin2    Lin3    -0.229
Kxr     Lx      Lin4    -0.138

.ends AQFP_RAM_CELL

.tran 0.05p 1800p 0 0.05p

.print i(Lin2.X1)
.print i(Id)
.print i(Iy)
.print i(Ix)
.print i(Iclk)
.print i(Lout)
* M test circuit

I1 0 1 pwl(0 0 10p 100u)
L1 1 0 2p
L2 2 0 2p
L3 2 0 0.2p
K1 L1 L2 0.2

.tran 0.25p 1600p 0 0.25p
.print i(L1) i(L2) i(L3)
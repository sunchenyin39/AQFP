* AQFP_BUFFER test circuit

Iin	    0	    1	    pwl(0 0 5p +20u)
Ixin	0	    2	    pwl(0 0 10p 0 20p 1.5m 1200p 1.5m 1220p 0)
X1      1       3       2       0       AQFP_BUFFER
Lout    3       0       6.8p

.subckt AQFP_BUFFER a q xin xout
.model jjmod jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param B1=0.5
.param B2=0.5
.param Lin=1.22p
.param Lx=5.19p
.param L1=1.42p
.param L2=1.42p
.param Lq=8.27p
.param Lout=28.4p
.param K1=-0.22
.param K2=-0.22
.param K3=+0.472
Lin     a       1       Lin
Lx      xin     xout    Lx
B1	    0	    2	    jjmod   area=B1
L1	    2	    1	    L1
L2	    1	    3	    L2
B2	    3	    0	    jjmod	area=B2
Lq	    1	    0	    Lq
Lout	q	    0	    Lout
K1	    Lx	    L1	    K1
K2	    Lx	    L2	    K2
K3	    Lq	    Lout	K3
.ends AQFP_BUFFER

.tran 0.25p 1600p 0 0.25p
.print i(Iin)
.print i(Ixin)
.print i(Lout)



